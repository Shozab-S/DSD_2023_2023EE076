`timescale 1ns / 1ps

module lab_4_tb;

    
    logic [1:0]a;
    logic [1:0]b;
    logic red, green, blue;
    
    
    lab_4 UUT (
        .a(a),
        .b(b),
        .red(red),
        .green(green),
        .blue(blue)
    );
    
    initial 
	begin
        
        a[0] = 0; a[1] = 0; b[0] = 0; b[1] = 0; 
		#10;
        a[0] = 0; a[1] = 0; b[0] = 1; b[1] = 0; 
		#10;
        a[0] = 0; a[1] = 0; b[0] = 0; b[1] = 1; 
		#10;
        a[0] = 0; a[1] = 0; b[0] = 1; b[1] = 1; 
		#10;
        a[0] = 1; a[1] = 0; b[0] = 0; b[1] = 0;
		#10;
        a[0] = 1; a[1] = 0; b[0] = 1; b[1] = 0; 
		#10;
        a[0] = 1; a[1] = 0; b[0] = 0; b[1] = 1; 
		#10;
        a[0] = 1; a[1] = 0; b[0] = 1; b[1] = 1; 
		#10;
        a[0] = 0; a[1] = 1; b[0] = 0; b[1] = 0; 
		#10;
        a[0] = 0; a[1] = 1; b[0] = 1; b[1] = 0;
		#10;
        a[0] = 0; a[1] = 1; b[0] = 0; b[1] = 1; 
		#10;
        a[0] = 0; a[1] = 1; b[0] = 1; b[1] = 1; 
		#10;
        a[0] = 1; a[1] = 1; b[0] = 0; b[1] = 0; 
		#10;
        a[0] = 1; a[1] = 1; b[0] = 1; b[1] = 0; 
		#10;
        a[0] = 1; a[1] = 1; b[0] = 0; b[1] = 1; 
		#10;
        a[0] = 1; a[1] = 1; b[0] = 1; b[1] = 1; 
        
        $stop;
    end
    
endmodule
